entity bcd is 
	port(a, b, c, d : in bit; s1, s2, s3, s4, s5, s6 : out bit);
end bcd;

architecture main of bcd is
	signal si1: bit;
	signal si2: bit;
	signal si3: bit;
	signal si4: bit;
	signal si5: bit;
	signal si6: bit;
begin
	-- Primeiro circuito que representa a saída s1
	
end architecture main;